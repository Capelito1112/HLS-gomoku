`timescale 1ns / 1ps

module pic_chess_piece(
    input wire can,
    input wire [31:0] y,
    output reg [28:0] ret
    );

    always @ (can or y)
        if (!can)
            ret = 23'b0;
        else
            case (y)
            32'd00: ret = 29'b00000000000111111100000000000;
            32'd01: ret = 29'b00000000111111111111100000000;
            32'd02: ret = 29'b00000011111111111111111000000;
            32'd03: ret = 29'b00000111111111111111111100000;
            32'd04: ret = 29'b00001111111111111111111110000;
            32'd05: ret = 29'b00011111111111111111111111000;
            32'd06: ret = 29'b00111111111111111111111111100;
            32'd07: ret = 29'b00111111111111111111111111100;
            32'd08: ret = 29'b01111111111111111111111111110;
            32'd09: ret = 29'b01111111111111111111111111110;
            32'd10: ret = 29'b01111111111111111111111111110;
            32'd11: ret = 29'b11111111111111111111111111111;
            32'd12: ret = 29'b11111111111111111111111111111;
            32'd13: ret = 29'b11111111111111111111111111111;
            32'd14: ret = 29'b11111111111111111111111111111;
            32'd15: ret = 29'b11111111111111111111111111111;
            32'd16: ret = 29'b11111111111111111111111111111;
            32'd17: ret = 29'b11111111111111111111111111111;
            32'd18: ret = 29'b01111111111111111111111111110;
            32'd19: ret = 29'b01111111111111111111111111110;
            32'd20: ret = 29'b01111111111111111111111111110;
            32'd21: ret = 29'b00111111111111111111111111100;
            32'd22: ret = 29'b00111111111111111111111111100;
            32'd23: ret = 29'b00011111111111111111111111000;
            32'd24: ret = 29'b00001111111111111111111110000;
            32'd25: ret = 29'b00000111111111111111111100000;
            32'd26: ret = 29'b00000011111111111111111000000;
            32'd27: ret = 29'b00000000111111111111100000000;
            32'd28: ret = 29'b00000000000111111100000000000;
            default: ret = 23'b0;
            endcase
    
endmodule

module pic_side_player(
    input wire can,
    input wire [31:0] y,
    output reg [71:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 72'b0;
        else
            case (y)
            32'd00: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 72'b001111111111111110000000011111000100000000001000010000010111111101111100;
            32'd04: ret = 72'b011111111111111111000000010000100100000000001000010000010100000001000010;
            32'd05: ret = 72'b011111111111111111000000010000010100000000010100001000100100000001000001;
            32'd06: ret = 72'b111111111111111111100000010000010100000000010100001000100100000001000001;
            32'd07: ret = 72'b111111111111111111100000010000010100000000010100000101000100000001000001;
            32'd08: ret = 72'b111111111111111111100000010000100100000000010100000101000100000001000010;
            32'd09: ret = 72'b111111111111111111100000011111000100000000100010000010000111111001111100;
            32'd10: ret = 72'b111111111111111111100000010000000100000000100010000010000100000001000100;
            32'd11: ret = 72'b111111111111111111100000010000000100000000100010000010000100000001000100;
            32'd12: ret = 72'b111111111111111111100000010000000100000000111110000010000100000001000010;
            32'd13: ret = 72'b011111111111111111000000010000000100000001000001000010000100000001000010;
            32'd14: ret = 72'b011111111111111111000000010000000100000001000001000010000100000001000001;
            32'd15: ret = 72'b001111111111111110000000010000000111111101000001000010000111111101000001;
            32'd16: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;
            default: ret = 72'b0;
            endcase
    
endmodule

module pic_side_ai(
    input wire can,
    input wire [31:0] y,
    output reg [71:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 72'b0;
        else
            case (y)
            32'd00: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 72'b001111111111111110000000000010000001110000000000000000000000000000000000;
            32'd04: ret = 72'b011111111111111111000000000010000000100000000000000000000000000000000000;
            32'd05: ret = 72'b011111111111111111000000000101000000100000000000000000000000000000000000;
            32'd06: ret = 72'b111111111111111111100000000101000000100000000000000000000000000000000000;
            32'd07: ret = 72'b111111111111111111100000000101000000100000000000000000000000000000000000;
            32'd08: ret = 72'b111111111111111111100000000101000000100000000000000000000000000000000000;
            32'd09: ret = 72'b111111111111111111100000001000100000100000000000000000000000000000000000;
            32'd10: ret = 72'b111111111111111111100000001000100000100000000000000000000000000000000000;
            32'd11: ret = 72'b111111111111111111100000001000100000100000000000000000000000000000000000;
            32'd12: ret = 72'b111111111111111111100000001111100000100000000000000000000000000000000000;
            32'd13: ret = 72'b011111111111111111000000010000010000100000000000000000000000000000000000;
            32'd14: ret = 72'b011111111111111111000000010000010000100000000000000000000000000000000000;
            32'd15: ret = 72'b001111111111111110000000010000010001110000000000000000000000000000000000;
            32'd16: ret = 72'b000111111111111100000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 72'b000011111111111000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 72'b000000111111100000000000000000000000000000000000000000000000000000000000;

            default: ret = 72'b0;
            endcase
    
endmodule

module pic_crt_ptr(
    input wire can,
    input wire [31:0] y,
    output reg [31:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 32'b0;
        else
            case (y)
            32'd00: ret = 32'b00000000000000000000000000000000;
            32'd01: ret = 32'b00000000000000000000000001000000;
            32'd02: ret = 32'b00000000000000000000000001100000;
            32'd03: ret = 32'b00000000000000000000000001110000;
            32'd04: ret = 32'b11111111111111111111111111111000;
            32'd05: ret = 32'b11111111111111111111111111111100;
            32'd06: ret = 32'b11111111111111111111111111111110;
            32'd07: ret = 32'b11111111111111111111111111111111;
            32'd08: ret = 32'b11111111111111111111111111111110;
            32'd09: ret = 32'b11111111111111111111111111111100;
            32'd10: ret = 32'b11111111111111111111111111111000;
            32'd11: ret = 32'b00000000000000000000000001110000;
            32'd12: ret = 32'b00000000000000000000000001100000;
            32'd13: ret = 32'b00000000000000000000000001000000;
            default: ret = 32'b0;
            endcase
    
endmodule


module pic_win(
    input wire can,
    input wire [31:0] y,
    output reg [85:0] ret
    );   
    
    always @ (can or y)
        if (!can)
            ret = 86'b0;
        else
            case (y)
                32'd00: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd01: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd02: ret = 86'b00000000000000000000000000000000000000000000000011100000000000000000000000000000000000;
                32'd03: ret = 86'b00000000000000000000000000000000000000000000000111111000000000000000000000000000000000;
                32'd04: ret = 86'b00000000000000000000000000000000000000000000011111111100000000000000000000000000000000;
                32'd05: ret = 86'b00000000000000000000000000000000000000000000011111111110000000000000000000000000000000;
                32'd06: ret = 86'b00000000000000000000000000000000000000000000011111111111000000000000000000000000000000;
                32'd07: ret = 86'b00000000000000000000000000000000000000000000011111111111000000000000000000000000000000;
                32'd08: ret = 86'b00000000000000000000001111000000000000000000011111111111000000000000000000000000000000;
                32'd09: ret = 86'b00000000000000000001111111110000000000000000011111111111111000000000000000000000000000;
                32'd10: ret = 86'b00000000000000000011111111111000000001000000001111111111111111000000000000000000000000;
                32'd11: ret = 86'b00000000111000000011111111111110000001110000000011111111111111110000000000000000000000;
                32'd12: ret = 86'b00000000111110000011111111111111000001111000000011111111111111111000000000000000000000;
                32'd13: ret = 86'b00000000111111000011111111111111000011111100000011111110001111111100000000000000000000;
                32'd14: ret = 86'b00000000111111110000000111111111000011111111111011111110000111111110000000000000000000;
                32'd15: ret = 86'b00000000111111111000000111111111000011111111111111111110001111111110000000000000000000;
                32'd16: ret = 86'b00000000111111111100000111111111000111111111111111111110011111111110000000000000000000;
                32'd17: ret = 86'b00000000011111111110000111111111000111111111111011111111111111111100000000000000000000;
                32'd18: ret = 86'b00000000011111111110000111111111000111111111110001111111111111110000000000000000000000;
                32'd19: ret = 86'b00000000011111111111000111111111000111111111100001111111111111110000000000000000000000;
                32'd20: ret = 86'b00000000011111111111000111111110000011111111100001111111111111000000000000000000000000;
                32'd21: ret = 86'b00000000001111111111000111111110000011111111111111111111111110000000000000000000000000;
                32'd22: ret = 86'b00000000001111111111111111111110000011111111111111111111111100000000000000000000000000;
                32'd23: ret = 86'b00000000001111111111111111111110000001111111111111111111111100000000000000000000000000;
                32'd24: ret = 86'b00000000001111111111111111111100000000001111111111111111111110000000000000000000000000;
                32'd25: ret = 86'b00000000001111111111111111111100000000001111111111111111111110000000000000000000000000;
                32'd26: ret = 86'b00000000001111111111111111111100000000001111111111111111111110000000000000000000000000;
                32'd27: ret = 86'b00000000001111111111111111111100000000001111111111111111111110000000000000000000000000;
                32'd28: ret = 86'b00000000001111111111111111111100000000000111111111111000111111111000000000000000000000;
                32'd29: ret = 86'b00000000001111111111110111111100000000000111111111111000011111111100000000000000000000;
                32'd30: ret = 86'b00000000011111111111001111111000000000000011111111111111111111111110000000000000000000;
                32'd31: ret = 86'b00000000011111111111001111111000000000001111111111111111111111111111000000000000000000;
                32'd32: ret = 86'b00000000011111111111001111111000000000111111111111111111111111111110000000000000000000;
                32'd33: ret = 86'b00000000011111111111011111111000000111111111111111111111111111111100000000000000000000;
                32'd34: ret = 86'b00000000011111111111111111111000011111111111111111111111111110000000000000000000000000;
                32'd35: ret = 86'b00000000011111111111111111111000111111111111111111111111100000000000000000000000000000;
                32'd36: ret = 86'b00000000011111111111111111111000111111111111111111111000000000000000000000000000000000;
                32'd37: ret = 86'b00000000011111111111111111111100111111111111111110111111111110000000000000000000000000;
                32'd38: ret = 86'b00000000111111111111111111111100111111111111111111111111111111111100000000000000000000;
                32'd39: ret = 86'b00000000111111111111111111111100111111111111111111111111101111111111000000000000000000;
                32'd40: ret = 86'b00000000111111111111111111111100011111111111111111111111110111111111110000000000000000;
                32'd41: ret = 86'b00000000111111111111111111111100000111111111110111111111111011111111111100000000000000;
                32'd42: ret = 86'b00000000111111111100001111111100001111111111100011111111111101111111111111000000000000;
                32'd43: ret = 86'b00000000111111111100001111111100001111111111000111111111111110111111111111100000000000;
                32'd44: ret = 86'b00000000111111111100001111111100111111111110001111111111111110011111111111110000000000;
                32'd45: ret = 86'b00000001111111111100001111111111111111111100111111111111111110011111111111111000000000;
                32'd46: ret = 86'b00000001111111111100001111111111111111111011111111111111111111101111111111111100000000;
                32'd47: ret = 86'b00000001111111111110001111111111111111111111111111111111111111110111111111111110000000;
                32'd48: ret = 86'b00000001111111111110000111111111111111111111111111111100011111111011111111111111000000;
                32'd49: ret = 86'b00000001111111111111000111111111111110111111111111111000111111111011111111111111000000;
                32'd50: ret = 86'b00000011111111111111100111111111110000111111111111110001111111111001111111111111000000;
                32'd51: ret = 86'b00000011111111111111100111111110000000000111111111100001111111111000001111111110000000;
                32'd52: ret = 86'b00000011111111101111111111111110000000001111111111000011111111111000000000000000000000;
                32'd53: ret = 86'b00000111111111001111111111111110000000011111111110000111111111111000000000000000000000;
                32'd54: ret = 86'b00000111111111000111111111111110000000111111111100001111111111111000000000000000000000;
                32'd55: ret = 86'b00000111111110000111111111111110000001111111111000011111111111110000000000000000000000;
                32'd56: ret = 86'b00001111111110000011111111111110000011111111110000111111111111110000000000000000000000;
                32'd57: ret = 86'b00001111111100000001111111111110000111111111100001111111111111100000000000000000000000;
                32'd58: ret = 86'b00011111111100000001111111111110001111111111100111111111111111100000000000000000000000;
                32'd59: ret = 86'b00011111111000000000111111111111011111111111111111111111111111000000000000000000000000;
                32'd60: ret = 86'b00111111111000000000111111111111000000001111111111111111111110000000000000000000000000;
                32'd61: ret = 86'b01111111110000000000011111111111000000001111111111111111111110000000000000000000000000;
                32'd62: ret = 86'b01111110000000000000011111111111000000000111111111111111111100000000000000000000000000;
                32'd63: ret = 86'b01111100000000000000001111111111000000000111111111111111111100000000000000000000000000;
                32'd64: ret = 86'b00000000000000000000000111111111000000000111111111111111110000000000000000000000000000;
                32'd65: ret = 86'b00000000000000000000000111111111000000000011111111111111100000000000000000000000000000;
                32'd66: ret = 86'b00000000000000000000000011111111000000000001111111111111000000000000000000000000000000;
                32'd67: ret = 86'b00000000000000000000000001111111000000000000111111111100000000000000000000000000000000;
                32'd68: ret = 86'b00000000000000000000000000011110000000000000011111111000000000000000000000000000000000;
                32'd69: ret = 86'b00000000000000000000000000000000000000000000011111100000000000000000000000000000000000;
                32'd70: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd71: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd72: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd73: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd74: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd75: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd76: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd77: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd78: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd79: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd80: ret = 86'b00000000000000000000000000000001111000000000000000000000000000000000000000000000000000;
                32'd81: ret = 86'b00000000000000000000000000000001111100000000000000000000000000000000000000000000000000;
                32'd82: ret = 86'b00000000000000000000000000000001111110000000000000000000000000000000000000000000000000;
                32'd83: ret = 86'b00000000000000000000000000000001111111000000000000000000000000000000000000000000000000;
                32'd84: ret = 86'b00000000000000000000000000000001111111100000000000000000000000000000000000000000000000;
                32'd85: ret = 86'b00000000000000000000000000000011111111100000000000000000000000000000000000000000000000;
                32'd86: ret = 86'b00000000000000000000000000000111111111100000000000000000000000000000000000000000000000;
                32'd87: ret = 86'b00000000000000000000000000001111111111101111111110000000000000000000000000000000000000;
                32'd88: ret = 86'b00000000000000000000000000011111111111111111111111000000000000000000000000000000000000;
                32'd89: ret = 86'b00000000000000000000000000111111111111111111111111100000000000000000000000000000000000;
                32'd90: ret = 86'b00000000000000000000000001111111111111111111111111110000000000000000000000000000000000;
                32'd91: ret = 86'b00000000000000000000001111111111111111111111111111111000000000000000000000000000000000;
                32'd92: ret = 86'b00000000000000000000001111111111111111111111111111111000000000000000000000000000000000;
                32'd93: ret = 86'b00000000000000000000011111111111111111111111111111111100000000000000000000000000000000;
                32'd94: ret = 86'b00000000000000000000111111111111111111111111111111111100000000000000000000000000000000;
                32'd95: ret = 86'b00000000000000000000111111111111111111111111111111111100000000000000000000000000000000;
                32'd96: ret = 86'b00000000000000000000111111111111110000111111111111111000000000000000000000000000000000;
                32'd97: ret = 86'b00000000000000000000111111111111000001111111111111110000000000000000000000000000000000;
                32'd98: ret = 86'b00000000000000000000111111111100000011111111111111100000000000000000000000000000000000;
                32'd99: ret = 86'b00000000000000000000111111110000000111111111111111000000000000000000000000000000000000;
                32'd100: ret = 86'b00000000000000000000111111100000001111111111111110000000000000000000000000000000000000;
                32'd101: ret = 86'b00000000000000000000011111000000111111111111111000000000000000000000000000000000000000;
                32'd102: ret = 86'b00000000000000000000001110000001111111111111110000000000000000000000000000000000000000;
                32'd103: ret = 86'b00000000000000000000000000000011111111111111100000000000000000000000000000000000000000;
                32'd104: ret = 86'b00000000000000000000000000000111111111111110000000000000000000000000000000000000000000;
                32'd105: ret = 86'b00000000000000000000000000111111111111111100000000000000000000000000000000000000000000;
                32'd106: ret = 86'b00000000000000000000000001111111111111111111111000000000000000000000000000000000000000;
                32'd107: ret = 86'b00000000000000000000000001111111111111111111111100000000000000000000000000000000000000;
                32'd108: ret = 86'b00000000000000000000000001111111111111111111111110000000000000000000000000000000000000;
                32'd109: ret = 86'b00000000000000000000000011111111111111111111111111000000000000000000000000000000000000;
                32'd110: ret = 86'b00000000000000000000000011111111111111111111111111100000000000000000000000000000000000;
                32'd111: ret = 86'b00000000000000000000000011111111111111111111111111100000000000000000000000000000000000;
                32'd112: ret = 86'b00000000000000000000000111111111000000000001111111100000000000000000000000000000000000;
                32'd113: ret = 86'b00000000000000000000000111111111111111110001111111100000000000000000000000000000000000;
                32'd114: ret = 86'b00000000000000000000001111111111111111111001111111100000000000000000000000000000000000;
                32'd115: ret = 86'b00000000000000000000001111111111111111111101111111100000000000000000000000000000000000;
                32'd116: ret = 86'b00000000000000000000001111111110011111111101111111110000000000000000000000000000000000;
                32'd117: ret = 86'b00000000000000000000011111111100011111111101111111110000000000000000000000000000000000;
                32'd118: ret = 86'b00000000000000000000011111111100011111111101111111110000000000000000000000000000000000;
                32'd119: ret = 86'b00000000000000000000111111111011111110000001111111110000000000000000000000000000000000;
                32'd120: ret = 86'b00000000000000000000111111111100000000000001111111110000000000000000000000000000000000;
                32'd121: ret = 86'b00000000000000000000111111111111111111100001111111110000000000000000000000000000000000;
                32'd122: ret = 86'b00000000000000000000111111111111111111110001111111110000000000000000000000000000000000;
                32'd123: ret = 86'b00000000000000000000111111111111111111110001111111110000000000000000000000000000000000;
                32'd124: ret = 86'b00000000000000000001111111110000011111110001111111111000000000000000000000000000000000;
                32'd125: ret = 86'b00000000000000000001111111110000111111110001111111111000000000000000000000000000000000;
                32'd126: ret = 86'b00000000000000000001111111100011111111100011111111111000000000000000000000000000000000;
                32'd127: ret = 86'b00000000000000000011111111100111111110011111111111111000000000000000000000000000000000;
                32'd128: ret = 86'b00000000000000000011111111101111000011111111111111111000000000000000000000000000000000;
                32'd129: ret = 86'b00000000000000000011111111111111111111111111111111111000000000000000000000000000000000;
                32'd130: ret = 86'b00000000000000000011111111111111111111111111111111111000000000000000000000000000000000;
                32'd131: ret = 86'b00000000000000000111111111111111111111111111111111111000000000000000000000000000000000;
                32'd132: ret = 86'b00000000000000000111111111111111111111111111111111111000000000000000000000000000000000;
                32'd133: ret = 86'b00000000000000000111111111111111111111111111111111111000000000000000000000000000000000;
                32'd134: ret = 86'b00000000000000000111111111111111111111111111111111111000000000000000000000000000000000;
                32'd135: ret = 86'b00000000000000000111111111111111111111111111111111111000000000000000000000000000000000;
                32'd136: ret = 86'b00000000000000000111111111111111111111111111111111110000000000000000000000000000000000;
                32'd137: ret = 86'b00000000000000000011111111111111111111100111111111000000000000000000000000000000000000;
                32'd138: ret = 86'b00000000000000000001111111111111111110000111111111110000000000000000000000000000000000;
                32'd139: ret = 86'b00000000000000000000011111111111111000000111111111111000000000000000000000000000000000;
                32'd140: ret = 86'b00000000000000001111111111111111110000000111111111111100000000000000000000000000000000;
                32'd141: ret = 86'b00000000000000011111111111111111000000000011111111111110000000000000000000000000000000;
                32'd142: ret = 86'b00000000000000111111111111111110000000000001111111111111000000000000000000000000000000;
                32'd143: ret = 86'b00000000000000111111111111111000000000000000111111111111100000000000000000000000000000;
                32'd144: ret = 86'b00000000000000111111111111110000000000000000011111111111110000000000000000000000000000;
                32'd145: ret = 86'b00000000000000111111111111100000000000000000001111111111110000000000000000000000000000;
                32'd146: ret = 86'b00000000000000111111111111000000000000000000001111111111110000000000000000000000000000;
                32'd147: ret = 86'b00000000000000111111111000000000000000000000000111111111110000000000000000000000000000;
                32'd148: ret = 86'b00000000000000111111110000000000000000000000000011111111110000000000000000000000000000;
                32'd149: ret = 86'b00000000000000111111100000000000000000000000000001111111100000000000000000000000000000;
                32'd150: ret = 86'b00000000000000011110000000000000000000000000000000111111100000000000000000000000000000;
                32'd151: ret = 86'b00000000000000000000000000000000000000000000000000011111000000000000000000000000000000;
                32'd152: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd153: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd154: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd155: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd156: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd157: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd158: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd159: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd160: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd161: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd162: ret = 86'b00000000000000000000000000000011111000000000000000000000000000000000000000000000000000;
                32'd163: ret = 86'b00000000000000000000000000001111111100000000000000000000000000000000000000000000000000;
                32'd164: ret = 86'b00000000000000000000000001111111111110000000000000000000000000000000000000000000000000;
                32'd165: ret = 86'b00000000000000000000000001111111111111000000000000000000000000000000000000000000000000;
                32'd166: ret = 86'b00000000000000000000000001111111111111110000000000000000000000000000000000000000000000;
                32'd167: ret = 86'b00000000000000000000000011111111111111111000000000000000000000000000000000000000000000;
                32'd168: ret = 86'b00000000000000000000000011111111100111111110000000000000000000000000000000000000000000;
                32'd169: ret = 86'b00000000000000000000000011111111000011111111100000000000000000000000000000000000000000;
                32'd170: ret = 86'b00000000000000000000000111111111000011111111110000000000000000000000000000000000000000;
                32'd171: ret = 86'b00000000000000000000000111111111000011111111111000000000000000000000000000000000000000;
                32'd172: ret = 86'b00000000000000000000001111111111000111111111111100000000000000000000000000000000000000;
                32'd173: ret = 86'b00000000000000000000001111111111001111111111111100000000000000000000000000000000000000;
                32'd174: ret = 86'b00000000000000000000001111111111111111111111111100000000000000000000000000000000000000;
                32'd175: ret = 86'b00000000000111100000011111111111111111111111111100000000000000000000000000000000000000;
                32'd176: ret = 86'b00000000000111111110011111111111111111111111111100000000000000000000000000000000000000;
                32'd177: ret = 86'b00000000000111111111111111111111111111111111111000000000000000000000000000000000000000;
                32'd178: ret = 86'b00000000000011111111111111111111111111111111100000000000000000000000000000000000000000;
                32'd179: ret = 86'b00000000000000111111111111111111111111111111000000000000000000000000000000000000000000;
                32'd180: ret = 86'b00000000000000011111111111111111111111111110000000000000000000000000000000000000000000;
                32'd181: ret = 86'b00000000000000001111111111111111111111110000000000000000000000000000000000000000000000;
                32'd182: ret = 86'b00000000000000000011111111111111111111000000000000000000000000000000000000000000000000;
                32'd183: ret = 86'b00000000000000000001111111111111110000000000000000000000000000000000000000000000000000;
                32'd184: ret = 86'b00000000000000000000111111111110000000011111100000000000000000000000000000000000000000;
                32'd185: ret = 86'b00000000000000000000111111111100000000111111110000000000000000000000000000000000000000;
                32'd186: ret = 86'b00000000000000000000111111111000000000011111111000000000000000000000000000000000000000;
                32'd187: ret = 86'b00000000000000000000111111111000000000001111111100000000000000000000000000000000000000;
                32'd188: ret = 86'b00000000000000000000111111111000000111111111111111000000000000000000000000000000000000;
                32'd189: ret = 86'b00000000000000000000111111111000111111111111111111110000000000000000000000000000000000;
                32'd190: ret = 86'b00000000000000000000111111111111111111111111111111111100000000000000000000000000000000;
                32'd191: ret = 86'b00000000000000000000111111111111111111111111111111111111000000000000000000000000000000;
                32'd192: ret = 86'b00000000000000000000111111111111111111111111111111111111100000000000000000000000000000;
                32'd193: ret = 86'b00000000000000000000111111111111111111111111111111111111110000000000000000000000000000;
                32'd194: ret = 86'b00000000000000000000111111111111111111001111111001111111111000000000000000000000000000;
                32'd195: ret = 86'b00000000000000000001111111111111111100011111111000011111111100000000000000000000000000;
                32'd196: ret = 86'b00000000000000000111111111111111110000011111110000011111111110000000000000000000000000;
                32'd197: ret = 86'b00000000000000001111111111111111000000111111110000001111111110000000000000000000000000;
                32'd198: ret = 86'b00000000000000011111111111111100000001111111110000000111111111000000000000000000000000;
                32'd199: ret = 86'b00000000000001111111111111111000000011111111100000000011111111100000000000000000000000;
                32'd200: ret = 86'b00000000000011111111111111111100000111111111100000000001111111110000000000000000000000;
                32'd201: ret = 86'b00000000000111111111111111111100001111111111000000000001111111111000000000000000000000;
                32'd202: ret = 86'b00000000001111111111111111111100011111111110000000000001111111111000000000000000000000;
                32'd203: ret = 86'b00000000011111111111111111111101111111111110000000000000111111111000000000000000000000;
                32'd204: ret = 86'b00000000111111111111101111111101111111111100000000000000111111111000000000000000000000;
                32'd205: ret = 86'b00000001111111111110001111111111111111111100000000000000111111111000000000000000000000;
                32'd206: ret = 86'b00000001111111111000001111111111111111111000000000000000111111111000000000000000000000;
                32'd207: ret = 86'b00000011111111100000000111111111111111100000000000000001111111111000000000000000000000;
                32'd208: ret = 86'b00000011111111000000000111111111111111000000000000000001111111111000000000000000000000;
                32'd209: ret = 86'b00000011111100000000000111111111111110000000000000000001111111111000000000000000000000;
                32'd210: ret = 86'b00000011111100000000011111111111111100000000000000000001111111111000000000000000000000;
                32'd211: ret = 86'b00000011111100000001111111111111110000000000000000000011111111111000000000000000000000;
                32'd212: ret = 86'b00000011111110000111111111111111110000000000000000000111111111111000000000000000000000;
                32'd213: ret = 86'b00000011111110011111111111111111110000000000000000001111111111110000000000000000000000;
                32'd214: ret = 86'b00000001111111111111111111111111110000000000000000011111111111100000000000000000000000;
                32'd215: ret = 86'b00000001111111111111111111111111110000000000000000111111111111100000000000000000000000;
                32'd216: ret = 86'b00000000111111111111111110000111110000000000000001111111111111000000000000000000000000;
                32'd217: ret = 86'b00000000011111111111111000000000000000000000000011111111111110000000000000000000000000;
                32'd218: ret = 86'b00000000011111111111000000000000000000000000000111111111111100000000000000000000000000;
                32'd219: ret = 86'b00000000000001110000000000000000000000000000011111111111111000000000000000000000000000;
                32'd220: ret = 86'b00000000000000000000000000000000000000000000111111111111110000000000000000000000000000;
                32'd221: ret = 86'b00000000000000000000000000000000000000000011111111111111000000000000000000000000000000;
                32'd222: ret = 86'b00000000000000000000000000000000000000001111111111111100000000000000000000000000000000;
                32'd223: ret = 86'b00000000000000000000000000000000000000111111111111110000000000000000000000000000000000;
                32'd224: ret = 86'b00000000000000000000000000000000000011111111111100000000000000000000000000000000000000;
                32'd225: ret = 86'b00000000000000000000000000000000000111111110000000000000000000000000000000000000000000;
                32'd226: ret = 86'b00000000000000000000000000000000000110000000000000000000000000000000000000000000000000;
                32'd227: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd228: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd229: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd230: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd231: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd232: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd233: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd234: ret = 86'b00000000000000000000000001100000000000000000000000000000000000000000000000000000000000;
                32'd235: ret = 86'b00000000000000000000000001110000000000000000000000000000000000000000000000000000000000;
                32'd236: ret = 86'b00000000000000000000000001111000000000000000000000000000000000000000000000000000000000;
                32'd237: ret = 86'b00000000000000000000000011111000000000000000000000000000000000000000000000000000000000;
                32'd238: ret = 86'b00000000000000000000000011111100000000011111000000000000000000000000000000000000000000;
                32'd239: ret = 86'b00000000000000000000000011111100000000011111100000000000000000000000000000000000000000;
                32'd240: ret = 86'b00000000000000000000000011111100000000011111110000000000000000000000000000000000000000;
                32'd241: ret = 86'b00000000000000000000000111111100000000001111111000000000000000000000000000000000000000;
                32'd242: ret = 86'b00000000000000000000000111111100000000001111111100000000000000000000000000000000000000;
                32'd243: ret = 86'b00000000000000000000001111111100000000001111111100000000000000000000000000000000000000;
                32'd244: ret = 86'b00000000000000000000001111111100000000001111111100000000000000000000000000000000000000;
                32'd245: ret = 86'b00000000000000000000011111111000000000001111111100000000000000000000000000000000000000;
                32'd246: ret = 86'b00000000000000000000011111111000000000001111111110000000000000000000000000000000000000;
                32'd247: ret = 86'b00000000000000000000011111111000000000001111111110000000000000000000000000000000000000;
                32'd248: ret = 86'b00000000000000000000111111111000000000001111111110000000000000000000000000000000000000;
                32'd249: ret = 86'b00000000000000000000111111111000000000001111111110000000000000000000000000000000000000;
                32'd250: ret = 86'b00000000000000000000111111110000000000001111111110000000000000000000000000000000000000;
                32'd251: ret = 86'b00000000000000000001111111110000000000001111111110000000000000000000000000000000000000;
                32'd252: ret = 86'b00000000000000000001111111110000000000001111111110000000000000000000000000000000000000;
                32'd253: ret = 86'b00000000000000000011111111100000000000001111111110000000000000000000000000000000000000;
                32'd254: ret = 86'b00000000000000000011111111100000000000001111111110000000000000000000000000000000000000;
                32'd255: ret = 86'b00000000000000000011111111100000000000001111111110000000000000000000000000000000000000;
                32'd256: ret = 86'b00000000000000000111111111000000000000001111111110000000000000000000000000000000000000;
                32'd257: ret = 86'b00000000000000000111111111000000000000001111111110000000000000000000000000000000000000;
                32'd258: ret = 86'b00000000000000000111111111100000000000001111111110000000000000000000000000000000000000;
                32'd259: ret = 86'b00000000000000000111111111100000000000001111111111000000000000000000000000000000000000;
                32'd260: ret = 86'b00000000000000001111111111100000000000001111111111000000000000000000000000000000000000;
                32'd261: ret = 86'b00000000000000001111111111100000000000001111111111000000000000000000000000000000000000;
                32'd262: ret = 86'b00000000000000001111111111100000000000001111111111000000000000000000000000000000000000;
                32'd263: ret = 86'b00000000000000001111111111100000000000001111111111000000000000000000000000000000000000;
                32'd264: ret = 86'b00000000000000001111111111100000000000001111111111000000000000000000000000000000000000;
                32'd265: ret = 86'b00000000000000001111111111100000000000001111111111000000000000000000000000000000000000;
                32'd266: ret = 86'b00000000000000001111111111100000000000001111111111000000000000000000000000000000000000;
                32'd267: ret = 86'b00000000000000001111111111000000000000001111111111000000000000000000000000000000000000;
                32'd268: ret = 86'b00000000000000001111111111000000000000001111111111000000000000000000000000000000000000;
                32'd269: ret = 86'b00000000000000001111111111000000000000001111111111000000000000000000000000000000000000;
                32'd270: ret = 86'b00000000000000000111111111000000000000001111111111000000000000000000000000000000000000;
                32'd271: ret = 86'b00000000000000000111111111000000000000001111111111000000000000000000000000000000000000;
                32'd272: ret = 86'b00000000000000000111111110000000000000001111111111000000000000000000000000000000000000;
                32'd273: ret = 86'b00000000000000000111111110000000000000001111111111000000000000000000000000000000000000;
                32'd274: ret = 86'b00000000000000000011111110000000000000001111111111000000000000000000000000000000000000;
                32'd275: ret = 86'b00000000000000000011111110000000000000001111111111000000000000000000000000000000000000;
                32'd276: ret = 86'b00000000000000000011111110000000000000001111111111000000000000000000000000000000000000;
                32'd277: ret = 86'b00000000000000000001111110000000000000001111111110000000000000000000000000000000000000;
                32'd278: ret = 86'b00000000000000000000111000000000000000001111111110000000000000000000000000000000000000;
                32'd279: ret = 86'b00000000000000000000000000000000000000001111111110000000000000000000000000000000000000;
                32'd280: ret = 86'b00000000000000000000000000000000000000011111111110000000000000000000000000000000000000;
                32'd281: ret = 86'b00000000000000000000000000000000000000011111111110000000000000000000000000000000000000;
                32'd282: ret = 86'b00000000000000000000000000000000000000011111111110000000000000000000000000000000000000;
                32'd283: ret = 86'b00000000000000000000000000000000000000011111111100000000000000000000000000000000000000;
                32'd284: ret = 86'b00000000000000000000000000000000000000011111111100000000000000000000000000000000000000;
                32'd285: ret = 86'b00000000000000000000000000000000000000011111111100000000000000000000000000000000000000;
                32'd286: ret = 86'b00000000000000000000000000000000000000011111111100000000000000000000000000000000000000;
                32'd287: ret = 86'b00000000000000000000000000000000000000011111111000000000000000000000000000000000000000;
                32'd288: ret = 86'b00000000000000000000000000000000000000111111111000000000000000000000000000000000000000;
                32'd289: ret = 86'b00000000000000000000000000000000000000111111111000000000000000000000000000000000000000;
                32'd290: ret = 86'b00000000000000000000000000000000000000111111111000000000000000000000000000000000000000;
                32'd291: ret = 86'b00000000000000000000000000000000000001111111110000000000000000000000000000000000000000;
                32'd292: ret = 86'b00000000000000000000000000000000000001111111110000000000000000000000000000000000000000;
                32'd293: ret = 86'b00000000000000000000000000000000000001111111110000000000000000000000000000000000000000;
                32'd294: ret = 86'b00000000000000000000000000000000000011111111100000000000000000000000000000000000000000;
                32'd295: ret = 86'b00000000000000000000000000000000000011111111100000000000000000000000000000000000000000;
                32'd296: ret = 86'b00000000000000000000000000000000000111111111100000000000000000000000000000000000000000;
                32'd297: ret = 86'b00000000000000000000000000000000000111111111000000000000000000000000000000000000000000;
                32'd298: ret = 86'b00000000000000000000000000000000001111111100000000000000000000000000000000000000000000;
                32'd299: ret = 86'b00000000000000000000000000000000011111111100000000000000000000000000000000000000000000;
                32'd300: ret = 86'b00000000000000000000000000000000011111111000000000000000000000000000000000000000000000;
                32'd301: ret = 86'b00000000000000000000000000000000111111110000000000000000000000000000000000000000000000;
                32'd302: ret = 86'b00000000000000000000000000000001111111100000000000000000000000000000000000000000000000;
                32'd303: ret = 86'b00000000000000000000000000000001111111000000000000000000000000000000000000000000000000;
                32'd304: ret = 86'b00000000000000000000000000000011111110000000000000000000000000000000000000000000000000;
                32'd305: ret = 86'b00000000000000000000000000000111111100000000000000000000000000000000000000000000000000;
                32'd306: ret = 86'b00000000000000000000000000000111111000000000000000000000000000000000000000000000000000;
                32'd307: ret = 86'b00000000000000000000000000000110000000000000000000000000000000000000000000000000000000;
                32'd308: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd309: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd310: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd311: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd312: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd313: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd314: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd315: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd316: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd317: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd318: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd319: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd320: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd321: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd322: ret = 86'b00000000000000000001111000000000000000000000000001111000000000000000000000000000000000;
                32'd323: ret = 86'b00000000000000000011111100000000000000000000000011111100000000000000000000000000000000;
                32'd324: ret = 86'b00000000000000000111111110000000000000000000000111111110000000000000000000000000000000;
                32'd325: ret = 86'b00000000000000000111111111000000000000000000000111111111000000000000000000000000000000;
                32'd326: ret = 86'b00000000000000001111111111000000000000000000001111111111000000000000000000000000000000;
                32'd327: ret = 86'b00000000000000001111111111000000000000000000001111111111000000000000000000000000000000;
                32'd328: ret = 86'b00000000000000001111111111100000000000000000001111111111100000000000000000000000000000;
                32'd329: ret = 86'b00000000000000001111111111100000000000000000001111111111100000000000000000000000000000;
                32'd330: ret = 86'b00000000000000001111111111100000000000000000001111111111100000000000000000000000000000;
                32'd331: ret = 86'b00000000000000001111111111100000000000000000001111111111100000000000000000000000000000;
                32'd332: ret = 86'b00000000000000001111111111100000000000000000001111111111100000000000000000000000000000;
                32'd333: ret = 86'b00000000000000001111111111100000000000000000001111111111100000000000000000000000000000;
                32'd334: ret = 86'b00000000000000001111111111000000000000000000001111111111000000000000000000000000000000;
                32'd335: ret = 86'b00000000000000001111111111000000000000000000001111111111000000000000000000000000000000;
                32'd336: ret = 86'b00000000000000001111111111000000000000000000001111111111000000000000000000000000000000;
                32'd337: ret = 86'b00000000000000001111111111000000000000000000001111111111000000000000000000000000000000;
                32'd338: ret = 86'b00000000000000001111111111000000000000000000001111111111000000000000000000000000000000;
                32'd339: ret = 86'b00000000000000001111111110000000000000000000001111111110000000000000000000000000000000;
                32'd340: ret = 86'b00000000000000001111111110000000000000000000001111111110000000000000000000000000000000;
                32'd341: ret = 86'b00000000000000001111111110000000000000000000001111111110000000000000000000000000000000;
                32'd342: ret = 86'b00000000000000001111111110000000000000000000001111111110000000000000000000000000000000;
                32'd343: ret = 86'b00000000000000011111111110000000000000000000011111111110000000000000000000000000000000;
                32'd344: ret = 86'b00000000000000011111111100000000000000000000011111111100000000000000000000000000000000;
                32'd345: ret = 86'b00000000000000011111111100000000000000000000011111111100000000000000000000000000000000;
                32'd346: ret = 86'b00000000000000011111111100000000000000000000011111111100000000000000000000000000000000;
                32'd347: ret = 86'b00000000000000011111111100000000000000000000011111111100000000000000000000000000000000;
                32'd348: ret = 86'b00000000000000011111111100000000000000000000011111111100000000000000000000000000000000;
                32'd349: ret = 86'b00000000000000111111111000000000000000000000111111111000000000000000000000000000000000;
                32'd350: ret = 86'b00000000000000111111111000000000000000000000111111111000000000000000000000000000000000;
                32'd351: ret = 86'b00000000000000111111111000000000000000000000111111111000000000000000000000000000000000;
                32'd352: ret = 86'b00000000000000111111111000000000000000000000111111111000000000000000000000000000000000;
                32'd353: ret = 86'b00000000000000111111111000000000000000000000111111110000000000000000000000000000000000;
                32'd354: ret = 86'b00000000000000111111111000000000000000000000111111110000000000000000000000000000000000;
                32'd355: ret = 86'b00000000000001111111111000000000000000000001111111110000000000000000000000000000000000;
                32'd356: ret = 86'b00000000000001111111110000000000000000000001111111110000000000000000000000000000000000;
                32'd357: ret = 86'b00000000000001111111110000000000000000000001111111100000000000000000000000000000000000;
                32'd358: ret = 86'b00000000000001111111110000000000000000000001111111100000000000000000000000000000000000;
                32'd359: ret = 86'b00000000000001111111100000000000000000000001111111100000000000000000000000000000000000;
                32'd360: ret = 86'b00000000000001111111100000000000000000000001111111000000000000000000000000000000000000;
                32'd361: ret = 86'b00000000000001111111100000000000000000000001111111000000000000000000000000000000000000;
                32'd362: ret = 86'b00000000000001111111000000000000000000000001111111000000000000000000000000000000000000;
                32'd363: ret = 86'b00000000000001111111000000000000000000000001111110000000000000000000000000000000000000;
                32'd364: ret = 86'b00000000000001111110000000000000000000000001111110000000000000000000000000000000000000;
                32'd365: ret = 86'b00000000000001111110000000000000000000000001111100000000000000000000000000000000000000;
                32'd366: ret = 86'b00000000000001111110000000000000000000000001111100000000000000000000000000000000000000;
                32'd367: ret = 86'b00000000000001111100000000000000000000000001111100000000000000000000000000000000000000;
                32'd368: ret = 86'b00000000000001111000000000000000000000000001110000000000000000000000000000000000000000;
                32'd369: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd370: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd371: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd372: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                32'd373: ret = 86'b00000000000011111000000000000000000000000011110000000000000000000000000000000000000000;
                32'd374: ret = 86'b00000000000011111000000000000000000000000011110000000000000000000000000000000000000000;
                32'd375: ret = 86'b00000000000111111000000000000000000000000111110000000000000000000000000000000000000000;
                32'd376: ret = 86'b00000000000111111100000000000000000000000111111000000000000000000000000000000000000000;
                32'd377: ret = 86'b00000000001111111100000000000000000000001111111000000000000000000000000000000000000000;
                32'd378: ret = 86'b00000000001111111100000000000000000000001111111000000000000000000000000000000000000000;
                32'd379: ret = 86'b00000000011111111100000000000000000000011111111000000000000000000000000000000000000000;
                32'd380: ret = 86'b00000000011111111100000000000000000000011111111000000000000000000000000000000000000000;
                32'd381: ret = 86'b00000000011111111100000000000000000000011111111000000000000000000000000000000000000000;
                32'd382: ret = 86'b00000000111111111100000000000000000000111111111000000000000000000000000000000000000000;
                32'd383: ret = 86'b00000000111111111100000000000000000000111111111000000000000000000000000000000000000000;
                32'd384: ret = 86'b00000000111111111100000000000000000000111111111000000000000000000000000000000000000000;
                32'd385: ret = 86'b00000000111111111100000000000000000000111111111000000000000000000000000000000000000000;
                32'd386: ret = 86'b00000000111111111100000000000000000000111111111000000000000000000000000000000000000000;
                32'd387: ret = 86'b00000000111111111100000000000000000000111111111000000000000000000000000000000000000000;
                32'd388: ret = 86'b00000000011111111100000000000000000000011111111000000000000000000000000000000000000000;
                32'd389: ret = 86'b00000000011111111000000000000000000000011111110000000000000000000000000000000000000000;
                32'd390: ret = 86'b00000000001111110000000000000000000000001111100000000000000000000000000000000000000000;
                32'd391: ret = 86'b00000000000111100000000000000000000000000111000000000000000000000000000000000000000000;
                32'd392: ret = 86'b00000000000110000000000000000000000000000100000000000000000000000000000000000000000000;
                32'd393: ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

            default: ret = 86'b0;
            endcase
    
endmodule

module pic_title(
    input wire can,
    input wire [31:0] y,
    output reg [85:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 86'b0;
        else
            case (y)
        32'd00:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd01:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd02:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd03:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd04:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd05:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd06:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd07:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd08:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd09:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd10:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd11:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd12:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd13:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd14:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd15:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd16:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd17:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd18:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd19:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd20:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd21:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd22:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd23:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd24:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd25:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd26:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd27:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd28:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd29:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd30:  ret = 86'b00000000000000000000000000000000000000000000000000000001111111111100000000000000000000;
        32'd31:  ret = 86'b00000000000000000000000000000000000000000000000001111111111111111110000000000000000000;
        32'd32:  ret = 86'b00000000000000000000000111000000000000000011111111111111111111111111000000000000000000;
        32'd33:  ret = 86'b00000000000000000000000111111111111111111111111111111111111111111111100000000000000000;
        32'd34:  ret = 86'b00000000000000000000000111111111111111111111111111111111111111111111110000000000000000;
        32'd35:  ret = 86'b00000000000000000000000011111111111111111111111111111111111111111111111000000000000000;
        32'd36:  ret = 86'b00000000000000000000000011111111111111111111111111111111111111111111111000000000000000;
        32'd37:  ret = 86'b00000000000000000000000001111111111111111111111111111111111111111111110000000000000000;
        32'd38:  ret = 86'b00000000000000000000000000111111111111111111111111111111111111111111110000000000000000;
        32'd39:  ret = 86'b00000000000000000000000000011111111111111111111111111111111111111110000000000000000000;
        32'd40:  ret = 86'b00000000000000000000000000000111111111111111111111111111111111000000000000000000000000;
        32'd41:  ret = 86'b00000000000000000000000000000000000111111111111111111100000000000000000000000000000000;
        32'd42:  ret = 86'b00000000000000000000000000000000000000000011111111111100000000000000000000000000000000;
        32'd43:  ret = 86'b00000000000000000000000000000000000000000011111111111100000000000000000000000000000000;
        32'd44:  ret = 86'b00000000000000000000000000000000000000000011111111111000000000000000000000000000000000;
        32'd45:  ret = 86'b00000000000000000000000000000000000000000111111111111000000000000000000000000000000000;
        32'd46:  ret = 86'b00000000000000000000000000000000000000000111111111110000000000000000000000000000000000;
        32'd47:  ret = 86'b00000000000000000000000000000000000000000111111111110000000000000000000000000000000000;
        32'd48:  ret = 86'b00000000000000000000000000000000000000001111111111110000000000000000000000000000000000;
        32'd49:  ret = 86'b00000000000000000000000000000000000000001111111111100000000000000000000000000000000000;
        32'd50:  ret = 86'b00000000000000000000000000000000000000011111111111100000000000000000000000000000000000;
        32'd51:  ret = 86'b00000000000000000000000000000000000000011111111111000000000000000000000000000000000000;
        32'd52:  ret = 86'b00000000000000000000000000000000000000111111111111000000000000000000000000000000000000;
        32'd53:  ret = 86'b00000000000000000000000000000000000000111111111111000000000000000000000000000000000000;
        32'd54:  ret = 86'b00000000000000000000000000000000000001111111111110000000000000000000000000000000000000;
        32'd55:  ret = 86'b00000000000000000000000000000000000011111111111111111100000000000000000000000000000000;
        32'd56:  ret = 86'b00000000000000000000000000000000001111111111111111111111111100000000000000000000000000;
        32'd57:  ret = 86'b00000000000000000000000000000011111111111111111111111111111111100000000000000000000000;
        32'd58:  ret = 86'b00000000000000000001111111111111111111111111111111111111111111110000000000000000000000;
        32'd59:  ret = 86'b00000000000000000001111111111111111111111111111111111111111111111000000000000000000000;
        32'd60:  ret = 86'b00000000000000000000111111111111111111111111111111111111111111111100000000000000000000;
        32'd61:  ret = 86'b00000000000000000000011111111111111111111111111111111111111111111110000000000000000000;
        32'd62:  ret = 86'b00000000000000000000001111111111111111111111111111111111111111111111000000000000000000;
        32'd63:  ret = 86'b00000000000000000000000111111111111111111111111111111111111111111111100000000000000000;
        32'd64:  ret = 86'b00000000000000000000000001111111111111111111110000000000111111111111100000000000000000;
        32'd65:  ret = 86'b00000000000000000000000000011111111111111111000000000000111111111111100000000000000000;
        32'd66:  ret = 86'b00000000000000000000000000001111111111111111000000000001111111111111100000000000000000;
        32'd67:  ret = 86'b00000000000000000000000000000011111111111110000000000001111111111111100000000000000000;
        32'd68:  ret = 86'b00000000000000000000000000000111111111111100000000000001111111111111000000000000000000;
        32'd69:  ret = 86'b00000000000000000000000000000111111111111000000000000001111111111111000000000000000000;
        32'd70:  ret = 86'b00000000000000000000000000001111111111111000000000000011111111111110000000000000000000;
        32'd71:  ret = 86'b00000000000000000000000000001111111111110000000000000011111111111110000000000000000000;
        32'd72:  ret = 86'b00000000000000000000000000011111111111110000000000000011111111111100000000000000000000;
        32'd73:  ret = 86'b00000000000000000000000000111111111111110000000000000111111111111100000000000000000000;
        32'd74:  ret = 86'b00000000000000000000000000111111111111100000000000000111111111111100000000000000000000;
        32'd75:  ret = 86'b00000000000000000000000001111111111111000000000000000111111111111000000000000000000000;
        32'd76:  ret = 86'b00000000000000000000000011111111111110000000000000001111111111111000000000000000000000;
        32'd77:  ret = 86'b00000000000000000000000111111111111100000000000000001111111111111000000000000000000000;
        32'd78:  ret = 86'b00000000000000000000011111111111111100000000000000011111111111110000000000000000000000;
        32'd79:  ret = 86'b00000000000000000000111111111111111000000000000000011111111111110000000000000000000000;
        32'd80:  ret = 86'b00000000000000000001111111111111110000000000000000111111111111100000000000000000000000;
        32'd81:  ret = 86'b00000000000000000001111111111111100000000000000001111111111111100000000000000000000000;
        32'd82:  ret = 86'b00000000000000000011111111111111111111111111111111111111111111111111111100000000000000;
        32'd83:  ret = 86'b00000000000000000011111111111111111111111111111111111111111111111111111111111110000000;
        32'd84:  ret = 86'b00000000000000111111111111111111111111111111111111111111111111111111111111111111000000;
        32'd85:  ret = 86'b00000000001111111111111111111111111111111111111111111111111111111111111111111111110000;
        32'd86:  ret = 86'b00000011111111111111111111111111111111111111111111111111111111111111111111111111111000;
        32'd87:  ret = 86'b00011111111111111111111111111111111111111111111111111111111111111111111111111111111000;
        32'd88:  ret = 86'b00011111111111111111111111111111111111111111111111111111111111111111111111111111111100;
        32'd89:  ret = 86'b00011111111111111111111111111111111111111111111111111111111111111111111111111111111100;
        32'd90:  ret = 86'b00001111111111111111111111111111111111111111111111111111111111111111111111111111111110;
        32'd91:  ret = 86'b00000111111111111111111111111111111110000000000000000000000111111111111111111111111110;
        32'd92:  ret = 86'b00000001111111111111111111110000000000000000000000000000000000000000011111111111111100;
        32'd93:  ret = 86'b00000000011111111110000000000000000000000000000000000000000000000000000000011111111100;
        32'd94:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd95:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd96:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd97:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd98:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd99:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd100:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd101:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd102:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd103:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd104:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd105:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd106:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd107:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd108:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd109:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd110:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd111:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd112:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd113:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd114:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd115:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd116:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd117:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd118:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd119:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd120:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd121:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd122:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd123:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd124:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd125:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd126:  ret = 86'b00000000000000000000000000000000000000000000000111111111111000000000000000000000000000;
        32'd127:  ret = 86'b00000000000000000000000000000000000000000001111111111111111111000000000000000000000000;
        32'd128:  ret = 86'b00000000000000000000000000000000000000000111111111111111111111100000000000000000000000;
        32'd129:  ret = 86'b00000000000000000000000000000000000000011111111111111111111111110000000000000000000000;
        32'd130:  ret = 86'b00000000000000000000000011100000000001111111111111111111111111111000000000000000000000;
        32'd131:  ret = 86'b00000000000000000000000011110000000111111111111111111111111111111100000000000000000000;
        32'd132:  ret = 86'b00000000000000000000000011111000001111111111111111111111111111111110000000000000000000;
        32'd133:  ret = 86'b00000000000000000000000011111110111111111111111111111111111111111111000000000000000000;
        32'd134:  ret = 86'b00000000000000000000000011111111111111111111111111111111111111111111000000000000000000;
        32'd135:  ret = 86'b00000000000000000000000011111111111111111100000000000000111111111111100000000000000000;
        32'd136:  ret = 86'b00000000000000000000000011111111111111000000000000000000111111111111110000000000000000;
        32'd137:  ret = 86'b00000000000000000000000011111111100000000000000000000000011111111111110000000000000000;
        32'd138:  ret = 86'b00000000000000000000000111111111000000000000000000000000011111111111110000000000000000;
        32'd139:  ret = 86'b00000000000000000000000111111110000000000000000000000000011111111111110000000000000000;
        32'd140:  ret = 86'b00000000000000000000000111111110000000000000000000000000011111111111110000000000000000;
        32'd141:  ret = 86'b00000000000000000000000111111110000000000000000000000000011111111111110000000000000000;
        32'd142:  ret = 86'b00000000000000000000000111111110000000011111111000000000011111111111110000000000000000;
        32'd143:  ret = 86'b00000000000000000000001111111110000111111111111111000000011111111111110000000000000000;
        32'd144:  ret = 86'b00000000000000000000001111111110011111111111111111100000011111111111110000000000000000;
        32'd145:  ret = 86'b00000000000000000000001111111111111111111111111111100000011111111111110000000000000000;
        32'd146:  ret = 86'b00000000000000000000001111111111111111111111111111110000011111111111110000000000000000;
        32'd147:  ret = 86'b00000000000000000000001111111111111111111111111111110000011111111111110000000000000000;
        32'd148:  ret = 86'b00000000000000000000001111111111111111111111111111110000011111111111110000000000000000;
        32'd149:  ret = 86'b00000000000000000000011111111111111111111111111111110000011111111111110000000000000000;
        32'd150:  ret = 86'b00000000000000000000011111111111111111111111111111110000011111111111110000000000000000;
        32'd151:  ret = 86'b00000000000000000000011111111111111111111111111111100000011111111111110000000000000000;
        32'd152:  ret = 86'b00000000000000000000011111111111111111111111111100000000011111111111110000000000000000;
        32'd153:  ret = 86'b00000000000000000000011111111111111111111111111100000000011111111111110000000000000000;
        32'd154:  ret = 86'b00000000000000000000011111111111110111111111100000000000011111111111110000000000000000;
        32'd155:  ret = 86'b00000000000000000000111111111110000111111111000000000000011111111111110000000000000000;
        32'd156:  ret = 86'b00000000000000000000111111111100001111111000000000000000011111111111110000000000000000;
        32'd157:  ret = 86'b00000000000000000000111111111100011111100000000000000000011111111111110000000000000000;
        32'd158:  ret = 86'b00000000000000000000111111111100111111000000000000000000011111111111110000000000000000;
        32'd159:  ret = 86'b00000000000000000000111111111101111100000111110000000000011111111111110000000000000000;
        32'd160:  ret = 86'b00000000000000000000111111111111111111111111111100000000011111111111110000000000000000;
        32'd161:  ret = 86'b00000000000000000000111111111111111111111111111110000000011111111111110000000000000000;
        32'd162:  ret = 86'b00000000000000000001111111111111111111111111111111000000011111111111110000000000000000;
        32'd163:  ret = 86'b00000000000000000001111111111111111111111111111111000000011111111111110000000000000000;
        32'd164:  ret = 86'b00000000000000000001111111111111111111111111111111000000011111111111110000000000000000;
        32'd165:  ret = 86'b00000000000000000001111111111111111111111111111111000000011111111111110000000000000000;
        32'd166:  ret = 86'b00000000000000000001111111111111111111111111111111000000011111111111110000000000000000;
        32'd167:  ret = 86'b00000000000000000011111111111111111111111111111110000000011111111111110000000000000000;
        32'd168:  ret = 86'b00000000000000000011111111111111111111111111111100000000011111111111110000000000000000;
        32'd169:  ret = 86'b00000000000000000011111111111111111111111111111000000000011111111111110000000000000000;
        32'd170:  ret = 86'b00000000000000000011111111111100000011111111100000000000011111111111110000000000000000;
        32'd171:  ret = 86'b00000000000000000011111111111000000011111111000000000000011111111111110000000000000000;
        32'd172:  ret = 86'b00000000000000000011111111111000000111111110000000000000011111111111110000000000000000;
        32'd173:  ret = 86'b00000000000000000011111111111000000111111100000000000000011111111111110000000000000000;
        32'd174:  ret = 86'b00000000000000000111111111111000001111111000000000000000011111111111110000000000000000;
        32'd175:  ret = 86'b00000000000000000111111111111000111111110000000000000000011111111111110000000000000000;
        32'd176:  ret = 86'b00000000000000000111111111111000111111100000000000000000011111111111110000000000000000;
        32'd177:  ret = 86'b00000000000000000111111111111001111111000000000000000000011111111111110000000000000000;
        32'd178:  ret = 86'b00000000000000000111111111111111111110000000000000000000011111111111110000000000000000;
        32'd179:  ret = 86'b00000000000000000111111111111111111100000000000000000000011111111111110000000000000000;
        32'd180:  ret = 86'b00000000000000000111111111111111111000000000000000000000011111111111110000000000000000;
        32'd181:  ret = 86'b00000000000000000111111111111111110000000000000000000000011111111111110000000000000000;
        32'd182:  ret = 86'b00000000000000000111111111111111111111111111111111111111111111111111110000000000000000;
        32'd183:  ret = 86'b00000000000000000111111111111111111111111111111111111111111111111111110000000000000000;
        32'd184:  ret = 86'b00000000000000000111111111111111111111111111111111111111111111111111110000000000000000;
        32'd185:  ret = 86'b00000000000000000111111111111111111111111111111111111111111111111111110000000000000000;
        32'd186:  ret = 86'b00000000000000000111111111111111111111111111111111111111111111111111110000000000000000;
        32'd187:  ret = 86'b00000000000000000011111111111111111111111111111111111111111111111111110000000000000000;
        32'd188:  ret = 86'b00000000000000000011111111111111111111111111111111111111111111111111110000000000000000;
        32'd189:  ret = 86'b00000000000000000001111111111111111111111111111111111111111111111111110000000000000000;
        32'd190:  ret = 86'b00000000000000000000111111111111111111111111111111111111111111111111110000000000000000;
        32'd191:  ret = 86'b00000000000000000000011111111111111111111111111111111111111111111111110000000000000000;
        32'd192:  ret = 86'b00000000000000000000000111111111111111111111111111111111111111111111110000000000000000;
        32'd193:  ret = 86'b00000000000000000000000001111111111111111111111111111111111111111111110000000000000000;
        32'd194:  ret = 86'b00000000000000000000000000000000000000000000000000000001111111111111110000000000000000;
        32'd195:  ret = 86'b00000000000000000000000000000000000000000000000000000001111111111111100000000000000000;
        32'd196:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111111000000000000000000;
        32'd197:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111110000000000000000000;
        32'd198:  ret = 86'b00000000000000000000000000000000000000000000000000000000011111111100000000000000000000;
        32'd199:  ret = 86'b00000000000000000000000000000000000000000000000000000000000111111000000000000000000000;
        32'd200:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd201:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd202:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd203:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd204:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd205:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd206:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd207:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd208:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd209:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd210:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd211:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd212:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd213:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd214:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd215:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd216:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd217:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd218:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd219:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd220:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd221:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd222:  ret = 86'b00000000000000000000000000000000000000000000000000000011100000000000000000000000000000;
        32'd223:  ret = 86'b00000000000000000000000000000011000000000000000001111111111100000000000000000000000000;
        32'd224:  ret = 86'b00000000000000000000000000001111000000000000111111111111111111000000000000000000000000;
        32'd225:  ret = 86'b00000000000000000000000000111111100000000111111111111111111111100000000000000000000000;
        32'd226:  ret = 86'b00000000000000000000000001111111100000111111111111111111111111111000000000000000000000;
        32'd227:  ret = 86'b00000000000000000000000011111111110111111111111110001111111111111100000000000000000000;
        32'd228:  ret = 86'b00000000000000000000000111111111111111111111100000001111111111111110000000000000000000;
        32'd229:  ret = 86'b00000000000000000000000111111111111111111110000000000111111111111111000000000000000000;
        32'd230:  ret = 86'b00000000000000000000001111111111111111111000000000001111111111111111000000000000000000;
        32'd231:  ret = 86'b00000000000000000000011111111111111111110000000000001111111111111111000000000000000000;
        32'd232:  ret = 86'b00000000000000000000011111111111111111100000000000011111111111111111000000000000000000;
        32'd233:  ret = 86'b00000000000000000000011111111111111111000000000000111111111111111111000000000000000000;
        32'd234:  ret = 86'b00000000000000000000011111111111111110000000000001111111111111111111000000000000000000;
        32'd235:  ret = 86'b00000000000000000000011111111111111100000000000011111111111111111110000000000000000000;
        32'd236:  ret = 86'b00000000000000000000011111111111111000000000001111111111111111111100000000000000000000;
        32'd237:  ret = 86'b00000000000000000000001111111111111000000000011111111111111111110000000000000000000000;
        32'd238:  ret = 86'b00000000000000000000001111111111111000000001111111111111111111000000000000000000000000;
        32'd239:  ret = 86'b00000000000000000000001111111111110000000011111111111111111110000000000000000000000000;
        32'd240:  ret = 86'b00000000000000000000000011111111110000001111111111111111111100000000000000000000000000;
        32'd241:  ret = 86'b00000000000000000000000011111111110000111111111111111111110000000000000000000000000000;
        32'd242:  ret = 86'b00000000000000000000000001111111100011111111111111111111111000000000000000000000000000;
        32'd243:  ret = 86'b00000000000000000000000000111111111111111111111111111111111100000000000000000000000000;
        32'd244:  ret = 86'b00000000000000000000000000000011111111111111111111111111111111000000000000000000000000;
        32'd245:  ret = 86'b00000000000000000000000000111111111111111111111111111111111111000000000000000000000000;
        32'd246:  ret = 86'b00000000000000000000001111111111111111111111111111111111111111000000000000000000000000;
        32'd247:  ret = 86'b00000000000000000000001111111111111111111111111111111111111111000000000000000000000000;
        32'd248:  ret = 86'b00000000000000000000001111111111111111111111111111111111111111000000000000000000000000;
        32'd249:  ret = 86'b00000000000000000000001111111111111111111111111111111111111110000000000000000000000000;
        32'd250:  ret = 86'b00000000000000000000000111111111111111111111111111111111111100000000000000000000000000;
        32'd251:  ret = 86'b00000000000000000000000011111111111111111111111111111111100000000000000000000000000000;
        32'd252:  ret = 86'b00000000000000000000000000111111111111111111111111111110000000000000000000000000000000;
        32'd253:  ret = 86'b00000000000000000000000000111111111111111111111111111100000000000000000000000000000000;
        32'd254:  ret = 86'b00000000000000000000000000011111111111111111111111111000000000000000000000000000000000;
        32'd255:  ret = 86'b00000000000000000000000000011111111111111111111111111000000000000000000000000000000000;
        32'd256:  ret = 86'b00000000000000000000000000011111111111111111111111111000000000000000000000000000000000;
        32'd257:  ret = 86'b00000000000000000000000000011111111111111111111111111000000000000000000000000000000000;
        32'd258:  ret = 86'b00000000000000000000000000011111111111110011111111111000000000000000000000000000000000;
        32'd259:  ret = 86'b00000000000000000000000000011111111111100011111111111000011111000000000000000000000000;
        32'd260:  ret = 86'b00000000000000000000000000011111111111100001111111111000111111110000000000000000000000;
        32'd261:  ret = 86'b00000000000000000000000000011111111111100001111111111001111111111000000000000000000000;
        32'd262:  ret = 86'b00000000000000000000000000011111111111100001111111111001111111111110000000000000000000;
        32'd263:  ret = 86'b00000000000000000000000000011111111111100001111111111001111111111111000000000000000000;
        32'd264:  ret = 86'b00000000000000000000000000011111111111100001111111111001111111111111100000000000000000;
        32'd265:  ret = 86'b00000000000000000000000000011111111111100001111111111000111111111111110000000000000000;
        32'd266:  ret = 86'b00000000000000001110000000011111111111100001111111111000001111111111111000000000000000;
        32'd267:  ret = 86'b00000000000000011111000000011111111111111001111111111000011111111111111000000000000000;
        32'd268:  ret = 86'b00000000000000111111110000011111111111111101111111111000011111111111111000000000000000;
        32'd269:  ret = 86'b00000000000000111111111000011111111111111101111111111000111111111111111000000000000000;
        32'd270:  ret = 86'b00000000000001111111111101111111111111111001111111111001111111111111110000000000000000;
        32'd271:  ret = 86'b00000000000001111111111111111111111111110001111111111011111111111111100000000000000000;
        32'd272:  ret = 86'b00000000000001111111111111111111111111100001111111111111111111111111000000000000000000;
        32'd273:  ret = 86'b00000000000011111111111111111111111111100001111111111111111111111100000000000000000000;
        32'd274:  ret = 86'b00000000000011111111111111111111111111100001111111111111111111111000000000000000000000;
        32'd275:  ret = 86'b00000000000011111111111111111111111111100001111111111111111111100000000000000000000000;
        32'd276:  ret = 86'b00000000000011111111111111111111111111100001111111111111111111000000000000000000000000;
        32'd277:  ret = 86'b00000000000011111111111111111111111111100001111111111111111110000000000000000000000000;
        32'd278:  ret = 86'b00000000000011111111111111011111111111100001111111111111110000000000000000000000000000;
        32'd279:  ret = 86'b00000000000011111111111100011111111111100001111111111111100000000000000000000000000000;
        32'd280:  ret = 86'b00000000000001111111111100011111111111100001111111111100000000000000000000000000000000;
        32'd281:  ret = 86'b00000000000000111111110000011111111111100001111111111000000000000000000000000000000000;
        32'd282:  ret = 86'b00000000000000011111100000011111111111100001111111111000000000000000000000000000000000;
        32'd283:  ret = 86'b00000000000000000000000000011111111111111001111111111000000000000000000000000000000000;
        32'd284:  ret = 86'b00000000000000000000000000011111111111111111111111111100000000000000000000000000000000;
        32'd285:  ret = 86'b00000000000000000000000000011111111111111111111111111100000000000000000000000000000000;
        32'd286:  ret = 86'b00000000000000000000000000011111111111111111111111111111111111111000000000000000000000;
        32'd287:  ret = 86'b00000000000000000000000000011111111111111111111111111111111111111111110000000000000000;
        32'd288:  ret = 86'b00000000000000000000000000011111111111111111111111111111111111111111111111100000000000;
        32'd289:  ret = 86'b00000000000000000000001111111111111111111111111111111111111111111111111111110000000000;
        32'd290:  ret = 86'b00000000000000000001111111111111111111111111111111111111111111111111111111111100000000;
        32'd291:  ret = 86'b00000000000000011111111111111111111111111111111111111111111111111111111111111110000000;
        32'd292:  ret = 86'b00000000000111111111111111111111111111111111111111111111111111111111111111111111000000;
        32'd293:  ret = 86'b00000011111111111111111111111111111111111111111111111111111111111111111111111111000000;
        32'd294:  ret = 86'b00111111111111111111111111111111111111111111111111111111111111111111111111111111100000;
        32'd295:  ret = 86'b00111111111111111111111111111111111111111111111111111111111111111111111111111111110000;
        32'd296:  ret = 86'b00111111111111111111111111111111110000000000000000000001111111111111111111111111110000;
        32'd297:  ret = 86'b00001111111111111111111111111110000000000000000000000000000000111111111111111111110000;
        32'd298:  ret = 86'b00000111111111111111111111110000000000000000000000000000000000000111111111111111110000;
        32'd299:  ret = 86'b00000011111111111111111100000000000000000000000000000000000000000001111111111111110000;
        32'd300:  ret = 86'b00000000111111111111110000000000000000000000000000000000000000000000000011111111000000;
        32'd301:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd302:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd303:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd304:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd305:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd306:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd307:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd308:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd309:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd310:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd311:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd312:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd313:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd314:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd315:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd316:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd317:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd318:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd319:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd320:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd321:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd322:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd323:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd324:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd325:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd326:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd327:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd328:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd329:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd330:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd331:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd332:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd333:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd334:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd335:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd336:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd337:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd338:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        32'd339:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000111111000000000;
        32'd340:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000111111111110000000;
        32'd341:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000011111111111111000000;
        32'd342:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000011111111111111100000;
        32'd343:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000011111111111111110000;
        32'd344:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000011111111111111110000;
        32'd345:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000001111111111111110000;
        32'd346:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000111111111111110000;
        32'd347:  ret = 86'b00000000000000000000000000000000000000000000000000000000000111111100001111111111110000;
        32'd348:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111111000001111111110000;
        32'd349:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111111111000000000000000;
        32'd350:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111111111100000000000000;
        32'd351:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111111111100000000000000;
        32'd352:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111111111110000000000000;
        32'd353:  ret = 86'b00000000000000000000000000000000000000000000000000000000011111111111111110000000000000;
        32'd354:  ret = 86'b00000000000000000000000000000000000000000000000000000000000111111111111110000000000000;
        32'd355:  ret = 86'b00000000000000000000000000000000000000000000000000000000000011111111111110000000000000;
        32'd356:  ret = 86'b00000000000000000000000000000000000000000000000000000000000001111111111110000000000000;
        32'd357:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000111111111100000000000000;
        32'd358:  ret = 86'b00000000000000000000000000000001111110000000000000000000000000001111100000000000000000;
        32'd359:  ret = 86'b00000000000000000000000000000111111111000000000000000000000000000000000000000000000000;
        32'd360:  ret = 86'b00000000000000000000000000011111111111100000000000000000000000000000000000000000000000;
        32'd361:  ret = 86'b00000000000000000000000011111111111111111000000000000000000000000000000000000000000000;
        32'd362:  ret = 86'b00000000000000000000001111111111111111111110000000000000000000000000000000000000000000;
        32'd363:  ret = 86'b00000000000011100000111111111111111111111111100000000000000000000000000000000000000000;
        32'd364:  ret = 86'b00000000001111100011111111111111111111111111111000000000000000000000000000000000000000;
        32'd365:  ret = 86'b00000000011111111111111111111111111111111111111100000000000000000000000000000000000000;
        32'd366:  ret = 86'b00000000011111111111111111111111111111111111111111000000000000000000000000000000000000;
        32'd367:  ret = 86'b00000000011111111111111111111111000011111111111111100000000000000000000000000000000000;
        32'd368:  ret = 86'b00000000011111111111111111111100000000111111111111111000000000000000000000000000000000;
        32'd369:  ret = 86'b00000000011111111111111111111000000000011111111111111100000000000000000000000000000000;
        32'd370:  ret = 86'b00000000011111111111111111100000000000000111111111111111000000000000000000000000000000;
        32'd371:  ret = 86'b00000000011111111111111110000000000000000011111111111111110000000000000000000000000000;
        32'd372:  ret = 86'b00000000001111111111111000000000000000000001111111111111111000000000000000000000000000;
        32'd373:  ret = 86'b00000000000111111111100000000000000000000000011111111111111110000000000000000000000000;
        32'd374:  ret = 86'b00000000000000000000000000000000000000000000001111111111111111000000000000000000000000;
        32'd375:  ret = 86'b00000000000000000000000000000000000000000000000111111111111111110000000000000000000000;
        32'd376:  ret = 86'b00000000000000000000000000000000000000000000000011111111111111111100000000000000000000;
        32'd377:  ret = 86'b00000000000000000000000000000000000000000000000001111111111111111111000000000000000000;
        32'd378:  ret = 86'b00000000000000000000000000000000000000000000000000011111111111111111100000000000000000;
        32'd379:  ret = 86'b00000000000000000000000000000000000000000000000000001111111111111111111100000000000000;
        32'd380:  ret = 86'b00000000000000000000000000000000000000000000000000000111111111111111111111000000000000;
        32'd381:  ret = 86'b00000000000000000000000000000000000000000000000000000001111111111111111111100000000000;
        32'd382:  ret = 86'b00000000000000000000000000000000000000000000000000000000111111111111111111111000000000;
        32'd383:  ret = 86'b00000000000000000000000000000000000000000000000000000000011111111111111111111100000000;
        32'd384:  ret = 86'b00000000000000000000000000000000000000000000000000000000000111111111111111111111000000;
        32'd385:  ret = 86'b00000000000000000000000000000000000000000000000000000000000001111111111111111111100000;
        32'd386:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000011111111111111111110000;
        32'd387:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000001111111111111111111000;
        32'd388:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000011111111111111111000;
        32'd389:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000011111111111111111000;
        32'd390:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000111111111111111000;
        32'd391:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111000;
        32'd392:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000111111111110000;
        32'd393:  ret = 86'b00000000000000000000000000000000000000000000000000000000000000000000000000111111100000;

            default: ret = 86'b0;
            endcase
    
endmodule

module pic_black_wins(
    input wire can,
    input wire [31:0] y,
    output reg [265:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 266'b0;
        else
            case (y)
            32'd00: ret = 266'b11111111111111111100000000000011111111000000000000000000000001111111111100000000000000000000011111100000000000000011111111000000000011111111110000000000000011111111000000011111111100000001111111100111111110000000111111100000000000111111100000000000000111110000000000;
            32'd01: ret = 266'b11111111111111111111100000000011111111000000000000000000000001111111111100000000000000000111111111111110000000000011111111000000000111111111100000000000000001111111000000011111111100000001111111000111111110000000111111110000000000111111100000000001111111111111000000;
            32'd02: ret = 266'b11111111111111111111110000000011111111000000000000000000000011111111111110000000000000011111111111111111100000000011111111000000001111111111000000000000000001111111000000011111111100000001111111000111111110000000111111110000000000111111100000000111111111111111110000;
            32'd03: ret = 266'b11111111111111111111111000000011111111000000000000000000000011111111111110000000000000111111111111111111110000000011111111000000011111111110000000000000000001111111100000111111111110000011111111000111111110000000111111111000000000111111100000001111111111111111111000;
            32'd04: ret = 266'b11111111111111111111111000000011111111000000000000000000000011111111111110000000000001111111111111111111111000000011111111000000111111111100000000000000000001111111100000111111111110000011111111000111111110000000111111111100000000111111100000011111111111111111111000;
            32'd05: ret = 266'b11111111111111111111111100000011111111000000000000000000000111111111111111000000000011111111111111111111111000000011111111000001111111111000000000000000000000111111100000111111111110000011111110000111111110000000111111111100000000111111100000011111111111111111111100;
            32'd06: ret = 266'b11111111000000011111111100000011111111000000000000000000000111111111111111000000000011111111100000011111111100000011111111000011111111110000000000000000000000111111100000111111111110000011111110000111111110000000111111111110000000111111100000111111111000001111111100;
            32'd07: ret = 266'b11111111000000001111111100000011111111000000000000000000000111111101111111000000000111111111000000001111111100000011111111000111111111100000000000000000000000111111110001111111111111000111111110000111111110000000111111111111000000111111100000111111110000000111111110;
            32'd08: ret = 266'b11111111000000001111111100000011111111000000000000000000000111111101111111000000000111111110000000000111111000000011111111001111111111000000000000000000000000111111110001111111111111000111111110000111111110000000111111111111000000111111100000111111110000000111000000;
            32'd09: ret = 266'b11111111000000001111111000000011111111000000000000000000001111111000111111100000000111111100000000000100000000000011111111011111111110000000000000000000000000111111110001111111111111000111111110000111111110000000111111111111100000111111100000111111111000000000000000;
            32'd10: ret = 266'b11111111000000011111111000000011111111000000000000000000001111111000111111100000000111111100000000000000000000000011111111111111111100000000000000000000000000011111110001111111111111000111111100000111111110000000111111111111110000111111100000011111111111100000000000;
            32'd11: ret = 266'b11111111111111111111110000000011111111000000000000000000001111111000111111100000001111111100000000000000000000000011111111111111111100000000000000000000000000011111110011111110111111100111111100000111111110000000111111111111110000111111100000011111111111111110000000;
            32'd12: ret = 266'b11111111111111111111100000000011111111000000000000000000011111111000011111110000001111111100000000000000000000000011111111111111111110000000000000000000000000011111111011111110111111101111111100000111111110000000111111101111111000111111100000001111111111111111100000;
            32'd13: ret = 266'b11111111111111111111000000000011111111000000000000000000011111110000011111110000001111111100000000000000000000000011111111111111111110000000000000000000000000011111111011111100011111101111111100000111111110000000111111101111111100111111100000000111111111111111111000;
            32'd14: ret = 266'b11111111111111111111110000000011111111000000000000000000011111110000011111110000001111111100000000000000000000000011111111111111111111000000000000000000000000001111111111111100011111111111111100000111111110000000111111100111111100111111100000000001111111111111111100;
            32'd15: ret = 266'b11111111111111111111111000000011111111000000000000000000111111110000001111111000001111111100000000000000000000000011111111111111111111100000000000000000000000001111111111111100011111111111111000000111111110000000111111100011111110111111100000000000001111111111111110;
            32'd16: ret = 266'b11111111111111111111111100000011111111000000000000000000111111111111111111111000001111111100000000000100000000000011111111111100111111100000000000000000000000001111111111111100011111111111111000000111111110000000111111100011111111111111100000000000000000111111111110;
            32'd17: ret = 266'b11111111000000001111111100000011111111000000000000000000111111111111111111111000000111111100000000000111100000000011111111111000011111110000000000000000000000001111111111111000001111111111111000000111111110000000111111100001111111111111100000000000000000000111111111;
            32'd18: ret = 266'b11111111000000000111111110000011111111000000000000000001111111111111111111111100000111111100000000000111111100000011111111110000011111110000000000000000000000001111111111111000001111111111111000000111111110000000111111100000111111111111100000000011100000000011111111;
            32'd19: ret = 266'b11111111000000000111111110000011111111000000000000000001111111111111111111111100000111111110000000001111111100000011111111100000001111111000000000000000000000000111111111111000001111111111110000000111111110000000111111100000011111111111100001111111100000000011111111;
            32'd20: ret = 266'b11111111000000000111111110000011111111000000000000000001111111111111111111111100000111111110000000011111111100000011111111000000001111111100000000000000000000000111111111110000000111111111110000000111111110000000111111100000011111111111100000111111110000000011111111;
            32'd21: ret = 266'b11111111000000001111111110000011111111111111111111000011111111111111111111111110000011111111000000111111111100000011111111000000000111111100000000000000000000000111111111110000000111111111110000000111111110000000111111100000001111111111100000111111111000000111111110;
            32'd22: ret = 266'b11111111111111111111111100000011111111111111111111000011111111111111111111111110000001111111111111111111111000000011111111000000000111111110000000000000000000000111111111110000000111111111110000000111111110000000111111100000000111111111100000111111111111111111111110;
            32'd23: ret = 266'b11111111111111111111111100000011111111111111111111000011111110000000000011111110000001111111111111111111111000000011111111000000000011111111000000000000000000000111111111110000000111111111110000000111111110000000111111100000000111111111100000011111111111111111111100;
            32'd24: ret = 266'b11111111111111111111111000000011111111111111111111000111111110000000000011111111000000111111111111111111110000000011111111000000000001111111000000000000000000000011111111100000000011111111100000000111111110000000111111100000000011111111100000001111111111111111111100;
            32'd25: ret = 266'b11111111111111111111111000000011111111111111111111000111111110000000000011111111000000011111111111111111100000000011111111000000000001111111100000000000000000000011111111100000000011111111100000000111111110000000111111100000000001111111100000000111111111111111110000;
            32'd26: ret = 266'b11111111111111111111100000000011111111111111111111000111111110000000000011111111000000000111111111111110000000000011111111000000000000111111110000000000000000000011111111100000000011111111100000000111111110000000111111100000000001111111100000000011111111111111100000;
            32'd27: ret = 266'b11111111111111110000000000000011111111111111111111001111111100000000000001111111100000000000011111100000000000000011111111000000000000111111110000000000000000000011111111100000000001111111100000000111111110000000111111100000000000111111100000000000000111111000000000;
            default: ret = 266'b0;
            endcase
    
endmodule

module pic_white_wins(
    input wire can,
    input wire [31:0] y,
    output reg [265:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 266'b0;
        else
            case (y)
            32'd00: ret = 266'b01111111100000001111111110000000111111110011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000001111111100000001111111110000000111111110011111111000000011111110000000000011111110000000000000011111000000000000;
            32'd01: ret = 266'b00111111100000001111111110000000111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111100000001111111110000000111111100011111111000000011111111000000000011111110000000000111111111111100000000;
            32'd02: ret = 266'b00111111100000001111111110000000111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111100000001111111110000000111111100011111111000000011111111000000000011111110000000011111111111111111000000;
            32'd03: ret = 266'b00111111110000011111111111000001111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111110000011111111111000001111111100011111111000000011111111100000000011111110000000111111111111111111100000;
            32'd04: ret = 266'b00111111110000011111111111000001111111100011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000111111110000011111111111000001111111100011111111000000011111111110000000011111110000001111111111111111111100000;
            32'd05: ret = 266'b00011111110000011111111111000001111111000011111111000000000111111110000000111111110000111111111111111111111111110000111111111111111111111100000000000000000011111110000011111111111000001111111000011111111000000011111111110000000011111110000001111111111111111111110000;
            32'd06: ret = 266'b00011111110000011111111111000001111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111110000011111111111000001111111000011111111000000011111111111000000011111110000011111111100000111111110000;
            32'd07: ret = 266'b00011111111000111111111111100011111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111111000111111111111100011111111000011111111000000011111111111100000011111110000011111111000000011111111000;
            32'd08: ret = 266'b00011111111000111111111111100011111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111111000111111111111100011111111000011111111000000011111111111100000011111110000011111111000000011100000000;
            32'd09: ret = 266'b00011111111000111111111111100011111111000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000011111111000111111111111100011111111000011111111000000011111111111110000011111110000011111111100000000000000000;
            32'd10: ret = 266'b00001111111000111111111111100011111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000001111111000111111111111100011111110000011111111000000011111111111111000011111110000001111111111110000000000000;
            32'd11: ret = 266'b00001111111001111111011111110011111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000001111111001111111011111110011111110000011111111000000011111111111111000011111110000001111111111111111000000000;
            32'd12: ret = 266'b00001111111101111111011111110111111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000001111111101111111011111110111111110000011111111000000011111110111111100011111110000000111111111111111110000000;
            32'd13: ret = 266'b00001111111101111110001111110111111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000001111111101111110001111110111111110000011111111000000011111110111111110011111110000000011111111111111111100000;
            32'd14: ret = 266'b00000111111111111110001111111111111110000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000000111111111111110001111111111111110000011111111000000011111110011111110011111110000000000111111111111111110000;
            32'd15: ret = 266'b00000111111111111110001111111111111100000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000000111111111111110001111111111111100000011111111000000011111110001111111011111110000000000000111111111111111000;
            32'd16: ret = 266'b00000111111111111110001111111111111100000011111111111111111111111110000000111111110000000000000111111110000000000000111111111111111111111000000000000000000000111111111111110001111111111111100000011111111000000011111110001111111111111110000000000000000011111111111000;
            32'd17: ret = 266'b00000111111111111100000111111111111100000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000111111111111100000111111111111100000011111111000000011111110000111111111111110000000000000000000011111111100;
            32'd18: ret = 266'b00000111111111111100000111111111111100000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000111111111111100000111111111111100000011111111000000011111110000011111111111110000000001110000000001111111100;
            32'd19: ret = 266'b00000011111111111100000111111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000011111111111100000111111111111000000011111111000000011111110000001111111111110000111111110000000001111111100;
            32'd20: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000011111111111000000011111111111000000011111111000000011111110000001111111111110000011111111000000001111111100;
            32'd21: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111110000000000000000000000000000000000011111111111000000011111111111000000011111111000000011111110000000111111111110000011111111100000011111111000;
            32'd22: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000011111111111000000011111111111000000011111111000000011111110000000011111111110000011111111111111111111111000;
            32'd23: ret = 266'b00000011111111111000000011111111111000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000011111111111000000011111111111000000011111111000000011111110000000011111111110000001111111111111111111110000;
            32'd24: ret = 266'b00000001111111110000000001111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000001111111110000000011111111000000011111110000000001111111110000000111111111111111111110000;
            32'd25: ret = 266'b00000001111111110000000001111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000001111111110000000011111111000000011111110000000000111111110000000011111111111111111000000;
            32'd26: ret = 266'b00000001111111110000000001111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000001111111110000000011111111000000011111110000000000111111110000000001111111111111110000000;
            32'd27: ret = 266'b00000001111111110000000000111111110000000011111111000000000111111110000000111111110000000000000111111110000000000000111111111111111111111100000000000000000000001111111110000000000111111110000000011111111000000011111110000000000011111110000000000000011111100000000000;
            default: ret = 266'b0;
            endcase
    
endmodule

module pic_res_draw(
    input wire can,
    input wire [31:0] y,
    output reg [265:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 266'b0;
        else
            case (y)
            32'd00: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000001111111111111111110000000000000000001111111111100000000001111111100000001111111110000000111111110000000000000000000000000000000000000000000000000000000000000000000000;
            32'd01: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000001111111111111111111110000000000000001111111111100000000000111111100000001111111110000000111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd02: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000001111111111111111111111100000000000011111111111110000000000111111100000001111111110000000111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd03: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111111111111111111110000000000011111111111110000000000111111110000011111111111000001111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd04: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111111111111111111110000000000011111111111110000000000111111110000011111111111000001111111100000000000000000000000000000000000000000000000000000000000000000000000;
            32'd05: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000001111111111111111111111110000000000111111111111111000000000011111110000011111111111000001111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd06: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000011111111100000001111111100000000111111111000000000111111111111111000000000011111110000011111111111000001111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd07: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000001111111110000001111111100000000011111111000000000111111101111111000000000011111111000111111111111100011111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd08: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000001111111100000000011111111000000000111111101111111000000000011111111000111111111111100011111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd09: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100000000011111111000000001111111000111111100000000011111111000111111111111100011111111000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd10: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100000000111111110000000001111111000111111100000000001111111000111111111111100011111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd11: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111111110000000001111111000111111100000000001111111001111111011111110011111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd12: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111111100000000011111111000011111110000000001111111101111111011111110111111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd13: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111111100000000011111110000011111110000000001111111101111110001111110111111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd14: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111110000000000011111110000011111110000000000111111111111110001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd15: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111000000000000111111110000001111111000000000111111111111110001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd16: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111111000001111111111111111111000000000000111111111111111111111000000000111111111111110001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd17: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100001111111100000000000111111111111111111111000000000111111111111100000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd18: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000011111110000001111111100000111111110000000001111111111111111111111100000000111111111111100000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd19: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000001111111100000011111111000000001111111111111111111111100000000011111111111100000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd20: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000001111111100000011111111000000001111111111111111111111100000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd21: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111100000001111111100000001111111100000001111111100000011111111111111111111111110000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd22: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000001111111100000001111111100000011111111111111111111111110000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd23: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111100000000111111110000011111110000000000011111110000000011111111111000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd24: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000001111111100000000011111111000111111110000000000011111111000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd25: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000001111111100000000011111111000111111110000000000011111111000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd26: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000001111111100000000001111111100111111110000000000011111111000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd27: ret = 266'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000001111111100000000001111111101111111100000000000001111111100000001111111110000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
            default: ret = 266'b0;
            endcase
    
endmodule

module pic_inst_draw(
    input wire can,
    input wire [31:0] y,
    output reg [604:0] ret
    );
    
    always @ (can or y)
        if (!can)
            ret = 605'b0;
        else
            case (y)
            32'd00: ret = 605'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd01: ret = 605'b01111111100000000000000000000000000000000000000000000000000000000000111110000001111111111101111100001111011111111111111011111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000001111000000111100011111110000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd02: ret = 605'b01111111110000000000000000000000000000000000000000000000000000000001111111100001111111111101111100001111011111111111111011111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111000000111100011111111000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd03: ret = 605'b01111111111000000000000000000000000000000000000000000000000000000011111111110001111111111101111100001111011111111111111011111111111011111111111000000000011100000000000000000000000000000000000111100000000000000000000000000011110000000000001111111111100000000000000000000000000000000000000000000000000001111000000111100011111111110000000000011100000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd04: ret = 605'b01111111111100000000000000000000000000000000000000000000000000000111111111111001111111111101111100001111011111111111111011111111111011111111111100000000011100000000000000000000000000000000000111100000000000000000000000000011110000000000001111111111110000000000000000000000000000000000000000000000000001111000000111100011111111111000000000011100000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd05: ret = 605'b01110000111110000000000000000000000000000000000000000000000000001111100011111001111111111101111100001111011111111111111011111111111011110001111100000000011100000000000000000000000000000000000111100000000000000000000000000011110000000000001111000011111000000000000000000000000000000000000000000000000001111000000111100011110011111100000000011100000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd06: ret = 605'b01110000011110000000000000000000000000000000000000000000000000011111000000110001110000000001111110001111000000111100000011100000000011110000111110000000011100000000000000000000000000000000000111100000000000000000000000000011110000000000001111000001111000000000000000000000000000000000000000000000000001111000000111100011110000111100000000011100000000000000000000000000000000000000000000000111000000000000000000000000000000111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd07: ret = 605'b01110000011110000000000000000000000000000000000000000000000000111111000000110001110000000001111110001111000000111100000011100000000011110000111110000000011100000000000000000000000000000000000111100000000000000000000000000011110000000000001111000001111000000000000000000000000000000000000000000000000001111000000111100011110000111100000000011100000000000000000000000000000000000000000000000111000000000000000000011110000000111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001110000000000000000000000000;
            32'd08: ret = 605'b01110000011110111100111000011111000000111111100001111100000000111110000000000001110000000001111110001111000000111100000011100000000011110000111110000001111111110000111110000000001111111000111111111100111111100000111001111111111111000000001111000001111011001111000011111100000111111000000111110000000001111000000111100011110000111100000001111111110000111111000000000011111100000001111100000111000000111111000000111111000111111110000000001111111110000111100001111110001111000001111000111111000011110111100000000111111000000110011111000000111110111100000000011111000000111111000001110000001111100000111001110;
            32'd09: ret = 605'b01110000011110111101111000111111100000111111110011111111000001111110000000000001110000000001111111001111000000111100000011100000000011110000111110000001111111110001111111100000001111111100111111111100111111110000111011111111111111000000001111000001111011011111000111111110001111111110001111111100000001111000000111100011110000111100000001111111110011111111100000000111111111000111111110000111000001111111100000111111110111111110000000001111111111000111100011111110000111100001111011111111100011110111100000001111111100000111111111100001111111111100000000111111110001111111100001110000111111111000111011110;
            32'd10: ret = 605'b01110000011110111111111001111111110001111111110111111111000001111100000000000001110000000001111111101111000000111100000011100000000011110000111100000001111111110011111111100000011111111100111111111100111111111000111111111111111111000000001111000001111011111111001111111110011111111110011111111100000001111000000111100011110000111100000001111111110111111111110000001111111111001111111111000111000011111111110001111111110111111110000000001111111111100111100011111111000111100011111011111111100011111111000000001111111110000111111111100011111111111100000001111111110011111111110001110001111111111100111111110;
            32'd11: ret = 605'b01110000011110111111111001111111110001111111110111111111000001111100000000000001110000000001111011101111000000111100000011100000000011110000111100000001111111110011111111100000011111111100111111111100111111111000111111111111111111000000001111000001111011111111001111111111011111111110011111111100000001111000000111100011110000111100000001111111110111111111111000011111111111001111111111000111000011111111110001111111110111111110000000001111111111110111100011111111000111100011111011111111100011111111000000001111111110000111111111110011111111111100000001111111110011111111110001110001111111111100111111110;
            32'd12: ret = 605'b01110000011110111111100011110001111001110000100111100010000001111100000000000001111111111001111011101111000000111100000011111111110011111111111100000000011100000111100011100000011100001000000111100000100001111000111111000011110000000000001111000001111011111000011110000111011110001100011100011000000001111000000111100011110001111100000000011100000111100001111000011111000010011111000111100111000111100001110011110001110000111000000000001111000011110111100010000111000011110011110111100001110011111110000000001100001111000111100011110111110001111100000011110001110111100001110001110001111000111100111111000;
            32'd13: ret = 605'b01111111111100111111000011100001111001110000000111100000000001111100000000000001111111111001111011111111000000111100000011111111110011111111111000000000011100000111000001110000011100000000000111100000000001111000111110000011110000000000001111111111110011110000011100000111011110000000011100000000000001111000000111100011111111111000000000011100000111000000111000011111000000011110000111100111000111000001110011100000000000111000000000001110000011110111100000000111000011110111110111000001110011111100000000000000001111000111000011110111100000111100000011110000000111000000111001110001110000011110111110000;
            32'd14: ret = 605'b01111111111100111110000011111111111001111110000111111000000001111100000000000001111111111001111011111111000000111100000011111111110011111111100000000000011100000111000001110000011111100000000111100000011111111000111100000011110000000000001111111111110011100000011111111111011111110000011111000000000001111000000111100011111111111000000000011100000111000000111000001111111000011111111111100111000111111111110011100000000000111000000000001110000001110111100001111111000001110111100111111111110011111100000000000011111111000111000001110111100000111100000011110000000111000000111001110001110000011110111100000;
            32'd15: ret = 605'b01111111111000111110000011111111111000111111100011111110000001111100000000000001110000000001111001111111000000111100000011100000000011111111110000000000011100000111000001110000001111111000000111100000111111111000111100000011110000000000001111111111000011100000011111111111001111111100001111111000000001111000000111100011111111100000000000011100000111000000111000000111111110011111111111100111000111111111110011100000000000111000000000001110000001110111100011111111000001111111100111111111110011111000000000001111111111000111000001110111100000111100000011110000000111000000111001110001110000011110111100000;
            32'd16: ret = 605'b01111111110000111110000011111111111000111111100011111110000001111100000000000001110000000001111001111111000000111100000011100000000011111111110000000000011100000111000001110000001111111000000111100000111111111000111100000011110000000000001111111111000011100000011111111110001111111100001111111000000001111000000111100011111111100000000000011100000111000000111000000111111110011111111111100111000111111111110011100000000000111000000000001110000001110111100011111111000001111111100111111111110011111000000000001111111111000111000001110111100000111100000011110000000111000000111001110001110000011110111100000;
            32'd17: ret = 605'b01110000000000111110000011111111111000011111110000111111000001111100000000000001110000000001111000111111000000111100000011100000000011110011111000000000011100000111000001110000000111111100000111100001111111111000111100000011110000000000001111000000000011100000011111111110000011111110000011111100000001111000000111100011110000000000000000011100000111000000111000000001111111011111111111100111000111111111110011100000000000111000000000001110000001110111100011111111000000111111000111111111110011111000000000011111111111000111000001110111100000111100000011110000000111000000111001110001110000011110111100000;
            32'd18: ret = 605'b01110000000000111110000011100000000000000111111000011111100001111110000000000001110000000001111000111111000000111100000011100000000011110001111000000000011100000111000001110000000001111110000111100001110001111000111100000011110000000000001111000000000011100000011100000000000000111111000011111110000001111000000111100011110000000000000000011100000111000000111000000000011111011110000000000111000111000000000011100000000000111000000000001110000011110111100011000111000000111111000111000000000011111000000000011110001111000111000001110111100000111100000011110000000111000000111001110001110000011110111100000;
            32'd19: ret = 605'b01110000000000111110000011100000010000000001111000000111100000111111000000110001110000000001111000011111000000111100000011100000000011110001111100000000011100000111000001110000000000011110000111100001110001111000111100000011110000000000001111000000000011100000011100000010000000001111000000111110000001111000000111100011110000000000000000011100000111000000111000000000000111011110000001000111000111000000010011100000000000111000000000001110000011110111100011000111000000011110000111000000000011111000000000011110001111000111000001110111100000111100000011110000000111000000111001110001110000011110111100000;
            32'd20: ret = 605'b01110000000000111110000011100000010000000001111000000111100000111111000000110001110000000001111000011111000000111100000011100000000011110001111100000000011100000111000001110000000000011110000111100001110001111000111100000011110000000000001111000000000011100000011100000111000000001111000000111110000001111000000111100011110000000000000000011100000111000000111000001000000111011110000001100111000111000000011011100000011000111000000000001110000011100111100011000111000000011110000111000000000011111000000000011110001111000111000001110111100000111100000011110000000111000000111001110001110000011110111100000;
            32'd21: ret = 605'b01110000000000111110000011110000111001100000111111000011100000011111100001111001110000000001111000011111000000111100000011100000000011110000111100000000011100000111100011100000011000001110000111100001110011111000111100000011110000000000001111000000000011100000011110000111011100001111011100011110000001111100001111100011110000000000000000011100000111100001111000001110000011011111000011100111000111100000111011110001111000111000000000001111111111100111100011000111000000011110000111100000110011111000000000011110001110000111000001110111110001111100000011110001110111100001110001110001111000111100111100000;
            32'd22: ret = 605'b01110000000000111110000001111111111001111111111111111111100000001111111111111001111111111101111000001111000000111100000011111111111011110000111110000000011111100011111111100000011111111110000111111001111111111000111100000011111110000111001111000000000011100000001111111111011111111111011111111110000001111111111111000011110000000000000000011111100111111111111000001111111111001111111111100111110011111111111001111111111000111110000000001111111111000111111011111111000000011100000011111111110011111000000000011111111110000111000001110011111111111100000001111111111011111111110001111101111111111100111100000;
            32'd23: ret = 605'b01110000000000111110000000111111110001111111110111111111000000000111111111111001111111111101111000001111000000111100000011111111111011110000011110000000011111110001111111100000011111111100000111111100111111111100111100000011111111001111101111000000000011100000001111111111011111111110011111111100000000111111111111000011110000000000000000011111110011111111110000001111111111000111111111000111110001111111110001111111110000111110000000001111111110000111111011111111100000111000000011111111100011111000000000001111111111000111000001110001111111111100000000111111110001111111100001111100111111111000111100000;
            32'd24: ret = 605'b01110000000000111110000000011111100000111111100011111110000000000011111111110001111111111101111000001111000000111100000011111111111011110000011111000000001111100001111111000000001111111000000011111000111110111100111100000001111110001111101111000000000011100000001111111110001111111100001111111000000000001111111110000011110000000000000000001111100001111111100000000111111110000011111110000111110001111111100000111111110000111110000000001110000000000111111001111111100111111000000001111111100011111000000000000111111111000111000001110000111111111100000000011111100001111111000001111100011111110000111100000;
            32'd25: ret = 605'b01110000000000111110000000011111100000111111100011111110000000000001111111100001111111111101111000001111000000111100000011111111111011110000011111000000001111100001111111000000001111111000000011111000111110111100111100000001111110000111101111000000000011100000000111111100001111111100001111111000000000000111111100000011110000000000000000001111100001111111000000000111111110000011111110000011110001111111100000111111100000111110000000001110000000000011111001111011100111111000000001111111100011111000000000000111111111000111000001110000111110111100000000011111100001111111000000111100011111110000111100000;
            32'd26: ret = 605'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd27: ret = 605'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd28: ret = 605'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            32'd29: ret = 605'b0;
            default: ret = 605'b0;
            endcase
endmodule
